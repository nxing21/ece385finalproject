//-------------------------------------------------------------------------
//    Ball.sv                                                            --
//    Viral Mehta                                                        --
//    Spring 2005                                                        --
//                                                                       --
//    Modified by Stephen Kempf     03-01-2006                           --
//                                  03-12-2007                           --
//    Translated by Joe Meng        07-07-2013                           --
//    Modified by Zuofu Cheng       08-19-2023                           --
//    Modified by Satvik Yellanki   12-17-2023                           --
//    Fall 2024 Distribution                                             --
//                                                                       --
//    For use with ECE 385 USB + HDMI Lab                                --
//    UIUC ECE Department                                                --
//-------------------------------------------------------------------------


module  ball 
( 
    input  logic        Reset, 
    input  logic        frame_clk,
    input  logic [7:0]  keycode,

    output logic [9:0]  BallX, 
    output logic [9:0]  BallY, 
    output logic [9:0]  BallS 
);
    

	 
    parameter [9:0] Ball_X_Center=320;  // Center position on the X axis
    parameter [9:0] Ball_Y_Center=24;  // Center position on the Y axis
    parameter [9:0] Ball_X_Min=224;       // Leftmost point on the X axis
    parameter [9:0] Ball_X_Max=420;     // Rightmost point on the X axis
    parameter [9:0] Ball_Y_Min=24;       // Topmost point on the Y axis
    parameter [9:0] Ball_Y_Max=460;     // Bottommost point on the Y axis
    parameter [9:0] Ball_X_Step=24;      // Step size on the X axis
    parameter [9:0] Ball_Y_Step=24;      // Step size on the Y axis

    logic [9:0] Ball_X_Motion;
    logic [9:0] Ball_X_Motion_next;
    logic [9:0] Ball_Y_Motion;
    logic [9:0] Ball_Y_Motion_next;

    logic [9:0] Ball_X_next;
    logic [9:0] Ball_Y_next;
    logic [7:0] prev_keycode;
    
    logic [7:0] timer;
    logic [7:0] downTick;
    
    logic alive;
    logic dummyAlive;

    always_comb begin
        Ball_Y_Motion_next = Ball_Y_Motion; // set default motion to be same as prev clock cycle 
        Ball_X_Motion_next = Ball_X_Motion;
        downTick = timer;
        dummyAlive = alive;

        //modify to control ball motion with the keycode
        if (keycode != 8'h00 && prev_keycode == 8'h00) begin
            if (keycode == 8'h1A) begin
                // Ball_Y_Motion_next = -10'd24;
                // Ball_X_Motion_next = 0;
            end else if (keycode == 8'h04 && dummyAlive) begin
                Ball_X_Motion_next = -10'd24;
                Ball_Y_Motion_next = 0;
            end else if (keycode == 8'h16) begin
                // Ball_Y_Motion_next = 10'd24;
                // Ball_X_Motion_next = 0;
            end else if (keycode == 8'h07 && dummyAlive) begin
                Ball_X_Motion_next = 10'd24;
                Ball_Y_Motion_next = 0;
            end
        end else begin
            Ball_X_Motion_next = 0;
            Ball_Y_Motion_next = 0;
        end
        
        if (downTick >= 50) begin
            if (BallY < Ball_Y_Max - BallS && dummyAlive) begin
                Ball_Y_Motion_next = 24;
            end else begin
                Ball_Y_Motion_next = 0;
            end
        end

//        if ( (BallY + BallS) >= Ball_Y_Max )  // Ball is at the bottom edge, BOUNCE!
//        begin
//            Ball_Y_Motion_next = (~ (Ball_Y_Step) + 1'b1);  // set to -1 via 2's complement.
//        end
//        else if ( (BallY - BallS) <= Ball_Y_Min )  // Ball is at the top edge, BOUNCE!
//        begin
//            Ball_Y_Motion_next = Ball_Y_Step;
//        end  
//       //fill in the rest of the motion equations here to bounce left and right
//        if ( (BallX + BallS) >= Ball_X_Max )
//        begin
//            Ball_X_Motion_next = (~ (Ball_X_Step) + 1'b1);
//        end
//        else if ( (BallX - BallS) <= Ball_X_Min )
//        begin
//            Ball_X_Motion_next = Ball_X_Step;
//        end
    end

    assign BallS = 24;  // default ball size
    assign Ball_X_next = (BallX + Ball_X_Motion_next);
    assign Ball_Y_next = (BallY + Ball_Y_Motion_next);
   
    always_ff @(posedge frame_clk) //make sure the frame clock is instantiated correctly
    begin: Move_Ball
        if (Reset)
        begin 
            Ball_Y_Motion <= 10'd0; //Ball_Y_Step;
			Ball_X_Motion <= 10'd0; //Ball_X_Step;
            
			BallY <= Ball_Y_Center;
			BallX <= Ball_X_Center;
			
			timer <= 0;
			downTick <= 0;
			alive <= 1;
			dummyAlive <= 1;
        end
        else 
        begin 
            
			Ball_Y_Motion <= Ball_Y_Motion_next; 
			Ball_X_Motion <= Ball_X_Motion_next; 
			
			if (!(Ball_Y_next > Ball_Y_Max || Ball_Y_next < Ball_Y_Min || Ball_X_next > Ball_X_Max || Ball_X_next < Ball_X_Min)) begin
                BallY <= Ball_Y_next;  // Update ball position
                BallX <= Ball_X_next;
            end
            
            prev_keycode <= keycode;
            timer <= timer + 1;
			
			if (timer >= 50) begin
			    timer <= 0;
			    
			    if (BallY > Ball_Y_Max - BallS) begin
			        alive <= 0;
			    end
			end
			
		end  
    end


    
      
endmodule
